package apb_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Define
    `include "apb_define.sv"
    `include "apb_master_transaction.sv"
    `include "apb_master_configuration.sv"

    // APB MASTER Components
    `include "apb_master_driver.sv"
    `include "apb_master_monitor.sv"
    `include "apb_master_sequencer.sv"
    `include "apb_master_coverage.sv"
    `include "apb_master_agent.sv"

endpackage : apb_pkg